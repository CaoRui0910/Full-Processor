module register32(q, d, clk, en, clr);
	input [31:0] d;
	input clk, en, clr;
	output [31:0] q;
	dffe1 dffe10(q[0], d[0], clk, en, clr);
	dffe1 dffe11(q[1], d[1], clk, en, clr);
	dffe1 dffe12(q[2], d[2], clk, en, clr);
	dffe1 dffe13(q[3], d[3], clk, en, clr);
	dffe1 dffe14(q[4], d[4], clk, en, clr);
	dffe1 dffe15(q[5], d[5], clk, en, clr);
	dffe1 dffe16(q[6], d[6], clk, en, clr);
	dffe1 dffe17(q[7], d[7], clk, en, clr);
	dffe1 dffe18(q[8], d[8], clk, en, clr);
	dffe1 dffe19(q[9], d[9], clk, en, clr);
	dffe1 dffe110(q[10], d[10], clk, en, clr);
	dffe1 dffe111(q[11], d[11], clk, en, clr);
	dffe1 dffe112(q[12], d[12], clk, en, clr);
	dffe1 dffe113(q[13], d[13], clk, en, clr);
	dffe1 dffe114(q[14], d[14], clk, en, clr);
	dffe1 dffe115(q[15], d[15], clk, en, clr);
	dffe1 dffe116(q[16], d[16], clk, en, clr);
	dffe1 dffe117(q[17], d[17], clk, en, clr);
	dffe1 dffe118(q[18], d[18], clk, en, clr);
	dffe1 dffe119(q[19], d[19], clk, en, clr);
	dffe1 dffe120(q[20], d[20], clk, en, clr);
	dffe1 dffe121(q[21], d[21], clk, en, clr);
	dffe1 dffe122(q[22], d[22], clk, en, clr);
	dffe1 dffe123(q[23], d[23], clk, en, clr);
	dffe1 dffe124(q[24], d[24], clk, en, clr);
	dffe1 dffe125(q[25], d[25], clk, en, clr);
	dffe1 dffe126(q[26], d[26], clk, en, clr);
	dffe1 dffe127(q[27], d[27], clk, en, clr);
	dffe1 dffe128(q[28], d[28], clk, en, clr);
	dffe1 dffe129(q[29], d[29], clk, en, clr);
	dffe1 dffe130(q[30], d[30], clk, en, clr);
	dffe1 dffe131(q[31], d[31], clk, en, clr);
endmodule
